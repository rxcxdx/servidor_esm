server {
  expires -1;
  root /home/rcd/apps/novo/dist;
}
